entity OR32 is
	port(
			a	:in bit_vector(31 downto 0);
			b	:in bit_vector(31 downto 0);
			output	:out bit_vector(31 downto 0)
		);
end OR32;
architecture test of OR32 is
begin
	output(0) <= a(0) or b(0);
	output(1) <= a(1) or b(1);
	output(2) <= a(2) or b(2);
	output(3) <= a(3) or b(3);
	output(4) <= a(4) or b(4);
	output(5) <= a(5) or b(5);
	output(6) <= a(6) or b(6);
	output(7) <= a(7) or b(7);
	output(8) <= a(8) or b(8);
	output(9) <= a(9) or b(9);
	output(10) <= a(10) or b(10);
	output(11) <= a(11) or b(11);
	output(12) <= a(12) or b(12);
	output(13) <= a(13) or b(13);
	output(14) <= a(14) or b(14);
	output(15) <= a(15) or b(15);
	output(16) <= a(16) or b(16);
	output(17) <= a(17) or b(17);
	output(18) <= a(18) or b(18);
	output(19) <= a(19) or b(19);
	output(20) <= a(20) or b(20);
	output(21) <= a(21) or b(21);
	output(22) <= a(22) or b(22);
	output(23) <= a(23) or b(23);
	output(24) <= a(24) or b(24);
	output(25) <= a(25) or b(25);
	output(26) <= a(26) or b(26);
	output(27) <= a(27) or b(27);
	output(28) <= a(28) or b(28);
	output(29) <= a(29) or b(29);
	output(30) <= a(30) or b(30);
	output(31) <= a(31) or b(31);
end test; 